module top (
    input logic clk,
    input logic rx,
    output logic tx
);

    assign tx = rx;

endmodule
